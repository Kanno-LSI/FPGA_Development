library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity autoencoder_tb is
end autoencoder_tb;

architecture Behavioral of autoencoder_tb is

component autoencoder
    Generic(
--        RAMaddressbit : integer := 13;
--        RAMaddressnum : integer := 8192;
        axi_bit : integer := 32;--PC�ʐM���̓��o�̓f�[�^��bit���B32bit�Œ�B
        data_dim : integer := 1024 ; --���́E�o�͑w�̑傫��(32�~32=1024)
        hide_dim : integer := 32 ; --�B��w�̑傫��
        data_bit : integer := 8 ; --���o�̓f�[�^��bit��
        weight_bit : integer := 16 ; --�d�݃f�[�^��bit��
        bias_bit : integer := 16 ;  --�o�C�A�X�f�[�^��bit��
        hide_bit : integer := 24 --�B��w�f�[�^��bit��
    );
    Port(
        CLK : in std_logic;
        X : in std_logic_vector(data_dim * data_bit -1 downto 0);
        ENCODE_START : in std_logic;
        Y : out std_logic_vector(data_dim * data_bit -1 downto 0);
        Y_ENABLE : out std_logic
    );
end component;

signal CLK_tb : std_LOGIC := '0';
signal ENCODE_START_tb : std_LOGIC := '0';
signal X_tb : std_logic_vector (8191 downto 0) := (others => '0');
signal Y_tb : std_logic_vector (8191 downto 0) := (others => '0');
signal Y_ENABLE_tb : std_LOGIC := '0';

begin
simulation_autoencoder : autoencoder port map(
    CLK => CLK_tb,
    ENCODE_START => ENCODE_START_tb,
    X  => X_tb,
    Y  => Y_tb,
    Y_ENABLE => Y_ENABLE_tb
);

process
begin
CLK_tb <= '0';
wait for 1 ns;
CLK_tb <= '1';
wait for 1 ns;
end process;

process
begin
ENCODE_START_tb <= '0';
wait for 3 ns;
wait for 100 ns;
ENCODE_START_tb <= '1';
wait for 2 ns;
ENCODE_START_tb <= '0';
wait for 40000 ns;
ENCODE_START_tb <= '1';
wait for 2 ns;
ENCODE_START_tb <= '0';
wait for 100000 ns;
end process;


process
begin
X_tb <=
--"01100100011000000110010101100001011000110110100001100100011010010111100001111101011100100111000101110111011111101000000110001000100100011001011110100001101010101011001010111011110000001100011011001101110101001110101011111000111101001110101111101110111011000110101001011111010111110101110101011111010111110110001101101110011111110111100101101101011010010110110001110010011110000111111010001000100011011001011010011101101000111010110010110101101110101100000111000101110100001101000011010100110110001101111011011000011000010101111101011010010110110101101001100000011011010111011110000000011111110110101101100001011000100110011001101010011101000111101110000001100010001001000010011010101000001010011010101011101011111011000110110110101110111100010011001011110100111100111001100000011001110110000001010101010101110110000101101010011100000111011001101110011011100110000101010011010111010110011001101111011101000111100001111110100001011000111110010100100110101001110110100010101001001010101010110011101110111100001111001010110001010101110101100010011001000100111101010111011000010110100001110000011010100110010101101010010110010100101001011110011011100111001101110100011101000111111110000111100001111000101110001101100100011001011110011101101001001010110010110111101111011100000010111010010101000110000001011101010100010101000001100101010111110110101101100000011001000110001001010101001111000101100001100101011010100111001101111110100000101000011001111110100000011000001010000110100011111001011010011111101010001011010010110101101110101011110101000011010011010100111101000011001111110100110001010001010110110101011001011111010101010100110001001011011000000110101001110010011101001000001001111101011101100111011101110011011110101000000110001001100011111001100010011110101001101010111110111110101101010011110001000110010000000011010100110100001101110011101100111111010000000100110101001001001111110100011101011001011011000110111001110101011101100111001001100111011010010111000101111010100000001000011110001111100101011001101110100011101010111011010110110000001101100011000100101111001011010010111000101111001100100011010100110110001110010011101000110010010011010101010001010101010110100110101101100100010111100101101001100001011100110111110010000010100001101000101110010000100110101010001010101001101011111010110000101000001010010010100100101000001010000010101000101110001100000010111100110001001100110010000000111010010001000100010001001001010100100101101001010010010100010110100001110100011111111000000110000010100010011000111110011100101000101010100110101011101001110001111000100011001001000010001000100011001001100010011000100011000100010001001100101100001010010011011000111011001111000011111101000011010001010100000101001010010100100101110101110011011101010111101010000111100010111001101010010111101001001010010110011011000010110001100100011111001000100010001000100010000111100001001000011001000111010001011000100011001010110010111100110011001110100011111000111111010000100100010001000011010001110101010001100010011011101000000110000111100011101001000010011011100101111000000100000011000001010001011100011100000110010001010100001111000111000010011000101001001000100001111000100110001010100010110000110000001101010011100000111110001111110100000001000001010001100100111101011000011010100111100101111110100010111001011001111100010110000001010100000111000010010001010000001111000110000010000100100110001010000010101100101001000101100001011000100000001001110010011000101001001100110011100100111100010000000100000101000100010001110100101101010100011000000110110001111111100010000101100101001011001001010010010100100100001000000010011100101001001010010010100100101010001011010010110000100100000110010001101000100010000110000010110100110100001101110011101000111011010000100100010101000110010010000100110101010100010111000110100001101101010011110101100000100001001010010010111000101101001011110011000000110001001100100011001100110101001101000011010000110001001010110010010100011010001001110011000000110011001100110010100100110010001111010100000101000100010001100100111101010110010111000101001001010111001110000001101100011111001011110011001000110011001101000011011100110110001101100011100000111010001111000011101000111001001110010011011100100111000111110001111100100101001011000010111100101100001110110100000001000001001111100011101100111111001100110011010000101110001001110010110100101110001100110011010000110110001110000011100000111001001110110011110000111111001111110100000001000000001111110011110100110000001011110011000100110011001100100010010100110000001110010011011000101111001010100011001100111101001100100100000100101000001100010011001000110000001100110011010100111000001110000011101000111011001111000011110101000000010000010100001001000010010000100100001101000101010001110100100101001001001110110011000000101011001010110011101100111001010000110100011001000101010011010011000100110101001101010011010100110110001110010011101100111100001111010011110100111110010000000100000101000100010001000100011001000110010001100100100001001001010011010100111101001110010011010100110001001000010010000011001101001001010011100100111101010011010000100011110100111101001111110100001101000011010000110100010001000100010001000100010101000110010011000101010001001001010011010101010001001011010010110100101001001100010011110101000101010010010100110101001001001100010000110100111101010011010110000110100100111100010001110100101101010001010101000101100001010101010100010101010001010010010101110101101001100101011000100100111101010000010111110101001101001110010011010100111001001110010100010101001101010100010100100100010001010010011000000110101001110001100000100100101001010111011000100111011001110100011100000111000001101100011011000110100001100101011010010110111101100101010110100101011001011011011000110101111101011000010100100101001001010011010101010101011001010110010101110101101101110100100001001000011110001110010101110101100001101011100010001001010010011010100101111001000010010000100011010111110001111111011110100111001001101001011001110110001001100111011010100110001101011110010111100101101001011000010101110101100001011001010110100111011010001001100011011000100001011111010111000110111010000001100110111001111110100001101001111010100110100001100110101010001010010101100001111000001001111101011100100111011101111001011110000111010101101110011101100110100001011011010110010101100001001000011010000111100110000011011111000110010101100110010111110111110110010001100101011001110010100010101010101010101110101100101100001010110010100011101000101001011010001101100101101001010110010010100001110111111001111010011111010110100001011110010110100101101001011111011010100111011101101100011010100110101001100001100000011000110010010101101000011010011010100101101010001010101110110000101101001011001010110111101011011010011010110010101101001010111010011001100011111000100010000001011101010110011001100001011000100101100001100011011010010110100101110110011100010110011101111010100010111001011110011100101001001010010110101010101011111011010110111011101111111011111110110011101110001011110111000001101101001010111010100110100110011001000101111011011011110110111001111001011011100110001101101001011011001000001001111011011110000111100110000101100101011001111110101000101011011011000110110000101101011011111111000100110001111011111110111011110000011100110010111111110000101011100010101110100111101000101101111100011110101000011110000001011110000110111001110000100011001000011110000110100000111000000010001101100101111010001010110000101101011011011010111001101111011100001011001010110011001100101111001010110100101100110011001010110001111100100110110100101000101000111110000111100101101001000101111110011101001000000010010010100011111001001110010110100110001001001010010101100111101010100010101011101100001011110011000011110010101100110111010010110011011101001111011001110110011101101011011101110101111100011010111110101001011001100010011111100101001000101010001000100011111001110010011001100101101001100110100010101001111001110010011010100111011010001110101011101101101011110111001100110100101101001011010111110100011101101111011111111001001110100111100111110101101100111011000000101011111010101110101110101000101010000010010100"
"10010010100100101001100110011101100110011001100110011101100110011001100110100000101001111010011110100111101001111010000010011101101000001010010010100111101001001010010010100100101000001010000010011101100100101001001010001011100001001000000001111100011100111000010010001110100101011001010110001110100100101001001010010010100100101001010110011101100111011001110110011001100101011001010110011001100111011001110110100000101001111010010010011101100111011001100110001011100001111000011101111100011100110111000001101010100001111000101110001110100011101000011110000111100010111000101110000111100010111000111010010010100011101000101110000100100010111000111010001110100100101001010110011101100101011000111010001110100011101000011101111001011111000111011001110011011011010110010110000000100001001000011110000111100001001000010010000000100000000111110010000000100001001000010010000100100000000111110001111100100000001000011110000111100100101001100110010010100001111000000010000100100000000111011001110000011100000110011101100101011001010111100101111100011111000111110001111001011110010111011001111001011110010111100101111001011100110111011001110110011110010111100101111100100000000111110010000111100010111000011110000000011111000111100101110110011100000110011101100111011000110101111001011110011100110111011001110011011100110111000001110000011011010111000001110000011100000110110101101101011100110111011001111001011101100111011001110110011100000111011010000100100000000111011001110110011100000111000001101010011000110101111001011100010110000101101001110000011100000110110101101101011001110110011101100111011010100110011101101010011001010110011101101010011100000111001101110000011011010110110101100111011100000111011001110110011011010111000001100111011010100110010101100000010111000101101001010111010101000110011101100111011001110110001101100000011000000101111001100011010111100110010101100000011000110110010101101010011010100110011101100101011000110110001101100101011010100110110101100111011001110110000001100011011000000101101001011010010110000101010101010100011000110110001101100000010111100101101001011010010110100101101001011010011000000101110001011100011000000110010101100111011000000110010101011100010110100101111001100011011001010110001101100011010111100101110001011010010110100101010101010101010101000101010001011110010111100101110001011000010101110101010101010100010101110101110001011110010101110101110001011110011000000110000001011100010111100101101001010111010111000101111001011110011000000110001101011100010110000101101001011000010101110101010101010100010100100101010101010101010101010101010001010100010100010101010101010111010110100101100001010101010110000101011101011000010110100101010101010101010101110101010001011000010110000101110001011100010111100101110001011000010101010101010101010101010101000101001001010010010100010101000101010001010100010101000101001111010100100101001001010100010101000101001001010101010101010101010001010101010100100101001001010100010100100101010001010111010110000101011101011110010111100101110001011000010101110101011101010111010101010101001001001111010011110100110101001101010011010100101101001111010011110100111101001101010100100101010001010010010011110100110101001101010011010100111101001111010100010101010001010010010101110101101001011010010110000101110001011100010110100101011101010101010101000100100001001000010010000100100001000101010000000100000001000101010000000100101101001101010011010100101101001011010010000100100001001000010010110100101101001111010011110101000101010101010101110101011101011000010111000101111001011100010111000101100001010100010000000100000001000000010000000100000001000000010000000011010101000000010000000100000001000000010000000100000001000000010000000100000001000101010001010100100001001101010011110101000101010001010100010101010101010111010110000101110001011100010110000101010000110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010101000000010000000100000001000000010000000100010101001011010011010100110101001111010100010101001001010101010110000101100001010111010110000011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010101000000010000000100000001000000010000000100000001000101010010000100101101001111010100100101010101010111010110000101100001011010001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010100000001000000010000000100000001000000010000000100000001000101010010110100111101010010010101000101011101011000010110000101010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101010000000100000001000000010000000100000001000000010000000100000001001000010010110100110101001111010100010101000101010010010011110011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010101000000010000000100000001000000010000000100000001000000010000000100000001000101010010000100100001001011010011010100110101001011001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010100000001000000010000000100000000110101001101010100000001000000010000000100000001000000010000000100000001000000010000000100000000110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010101000000010000000100000001000000010000000100000001000000010000000011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101010000000100000001000000010000000100000000110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101010000000100000000110101001101010011010100110101001101010011010100110101001101010011010100110101001101010011010100110101"
;
wait for 5 ns;
end process;




end Behavioral;
